magic
tech sky130A
timestamp 1628866758
<< error_p >>
rect -33 700 233 733
rect -33 0 0 700
rect 200 0 233 700
rect -33 -33 233 0
<< mvnsubdiff >>
rect 0 690 200 700
rect 0 10 10 690
rect 190 10 200 690
rect 0 0 200 10
<< mvnsubdiffcont >>
rect 10 10 190 690
<< locali >>
rect 0 690 200 700
rect 0 10 10 690
rect 190 10 200 690
rect 0 0 200 10
<< viali >>
rect 10 10 190 690
<< metal1 >>
rect 0 690 200 700
rect 0 10 10 690
rect 190 10 200 690
rect 0 0 200 10
<< via1 >>
rect 10 10 190 690
<< metal2 >>
rect 0 690 200 700
rect 0 10 10 690
rect 190 10 200 690
rect 0 0 200 10
<< via2 >>
rect 10 10 190 690
<< metal3 >>
rect 0 690 200 700
rect 0 10 10 690
rect 190 10 200 690
rect 0 0 200 10
<< end >>
