magic
tech sky130A
timestamp 1628793935
<< mvnmos >>
rect 0 0 100 2000
<< mvndiff >>
rect -52 0 0 2000
rect 100 0 150 2000
<< poly >>
rect 0 2000 100 2050
rect 0 -50 100 0
<< end >>
