magic
tech sky130A
timestamp 1628867017
<< mvpsubdiff >>
rect 0 680 200 700
rect 0 20 20 680
rect 180 20 200 680
rect 0 0 200 20
<< mvpsubdiffcont >>
rect 20 20 180 680
<< locali >>
rect 0 680 200 700
rect 0 20 20 680
rect 180 20 200 680
rect 0 0 200 20
<< viali >>
rect 20 20 180 680
<< metal1 >>
rect 0 680 200 700
rect 0 20 20 680
rect 180 20 200 680
rect 0 0 200 20
<< end >>
