magic
tech sky130A
timestamp 1628793262
<< mvnmos >>
rect 0 0 500 2000
<< mvndiff >>
rect -100 0 0 2000
rect 500 0 600 2000
<< poly >>
rect 0 2000 500 2050
rect 0 -50 500 0
<< end >>
