magic
tech sky130A
timestamp 1628865753
<< error_p >>
rect -23 90 123 123
rect 4 86 123 90
rect 4 84 14 86
rect 10 14 14 84
rect 86 14 123 86
rect 10 10 123 14
rect 84 4 123 10
rect 90 -23 123 4
<< mvpdiffc >>
rect 10 10 90 90
<< locali >>
rect 0 90 100 100
rect 0 10 10 90
rect 90 10 100 90
rect 0 0 100 10
<< viali >>
rect 10 10 90 90
<< metal1 >>
rect 0 90 100 100
rect 0 10 10 90
rect 90 10 100 90
rect 0 0 100 10
<< end >>
