*ANALOG BANDGAP REFERENCE CIRCUIT  

*STARTUP_CHECK

.options savecurrents
.lib "sky130_fd_pr/models/sky130.lib.spice" tt
.include "sky130_fd_pr/models/sky130_fd_pr__model__pnp.model.spice"

*BGR CIRCUIT

.option scale=0.005u

X0 F VREF VSSA sky130_fd_pr__res_xhigh_po w=70 l=9604
X3 E J VSSA sky130_fd_pr__res_xhigh_po w=70 l=1079
X7 K VDDB VSSA sky130_fd_pr__res_xhigh_po w=70 l=6998

X1 sky130_fd_pr__pnp_05v5_W3p40L3p40_0/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_0/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X2 sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X4 sky130_fd_pr__pnp_05v5_W3p40L3p40_3/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_3/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X5 sky130_fd_pr__pnp_05v5_W3p40L3p40_2/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_2/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X6 sky130_fd_pr__pnp_05v5_W3p40L3p40_4/c_153_607# VSSA I sky130_fd_pr__pnp_05v5_W3p40L3p40_4/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X8 sky130_fd_pr__pnp_05v5_W3p40L3p40_5/c_153_607# VSSA F sky130_fd_pr__pnp_05v5_W3p40L3p40_5/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X9 sky130_fd_pr__pnp_05v5_W3p40L3p40_6/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_6/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X10 sky130_fd_pr__pnp_05v5_W3p40L3p40_7/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_7/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X11 sky130_fd_pr__pnp_05v5_W3p40L3p40_8/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_8/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X13 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1

X12 B En I VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=113 ps=0 w=4000 l=1000
X14 D A C VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X15 A A B VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X16 J En D VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=-1 pd=-1 as=0 ps=0 w=4000 l=1000
X17 H En VREF VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X18 C G VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X19 G En K VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X20 G A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=200
X21 A C VDDB VDDB sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X22 C C VDDB VDDB sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X23 H C VDDB VDDB sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000

C0 K G 0.25fF
C1 K VREF 0.27fF
C2 G A 0.12fF
C3 C VREF 0.55fF
C4 A VREF 0.28fF
C5 C En 0.61fF
C6 En A 0.53fF
C7 VDDB C 0.09fF
C8 VDDB A 0.10fF
C9 I A 0.12fF
C10 I J 0.28fF
C11 C A 0.67fF
C12 G En 0.65fF
C13 En VREF 0.22fF
C14 H VDDB 0.04fF
C15 VDDB VSSA 82.44fF
C16 E VSSA 4.86fF

R3 GND VREF 100MEG

VSS VSSA GND DC 0V
VD En GND DC 3.3V

VDD VDDB GND pulse(0V 3.3V 100u 100u 0 0.5 1 0)


.tran 1u 900u

.control

run

plot V(EN)
plot -I(Vdd)

.endc

.end


