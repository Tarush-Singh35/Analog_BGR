magic
tech sky130A
timestamp 1628792784
<< nwell >>
rect -251 -151 750 2150
<< mvpmos >>
rect 0 0 500 2001
<< mvpdiff >>
rect -100 0 0 2001
rect 500 0 600 2001
<< poly >>
rect 0 2001 500 2025
rect 0 -25 500 0
<< end >>
